/********************************************************************
 *                TEST BENCH FOR PROTECTION CELLS                   *
 ********************************************************************
 * Laboratory    : Robotics and Embedded System Technology
 * Engineer      : Hanjara Cahya Adhyatma
 * Create Date   : 12/05/2017
 * Project Name  : FINAL PROJECT
 * Target Devices: TEST BENCH SIM PROTECTION AND FPGA
 * Tool versions : VERILOG 2001 RUN ON ICARUS 10
 * Description   :　日本へかえりますために。。。
 * Dependencies  :　いない
 * Revision      :　今から
 * Additional Comments:　いない
 ********************************************************************
 *                       INCLUDE MODULES                            *
 *******************************************************************/
`include "../module/top.v"
/********************************************************************
 *                        IO DEFINITIONS                            *
 *******************************************************************/
module protection_sim;
	reg [3:0] a, b;
	wire [7:0] c;
/********************************************************************
 *                         DUMPER MONITOR                           *
 *******************************************************************/
	initial
	begin
		$dumpfile("vcd");
		$dumpvars(0, tops);
		$monitor($time, " A=%d b=%d a*b=%d",a,b,c);
	end
/********************************************************************
 *                            CLOCKING                              *
 *******************************************************************
	initial
	begin
		CLK  = 1'b1;
		forever #5 CLK = ~CLK;
	end
 ********************************************************************
 *                              RESET                               *
 *******************************************************************
	initial 
	begin
		RST = 1'b1;
		#5 RST = 1'b0;
	end
 ********************************************************************
 *                         DATAS INJECTION                          *
 *******************************************************************/
	initial
	begin
		a = 3'b000;
		#2 a = 3'b001;
		#2 a = 3'b010;
		#2 a = 3'b011;
		#2 a = 3'b100;

	end

	initial
	begin
		b = 3'b000;
		#2 b = 3'b010;
		#2 b = 3'b010;
		#2 b = 3'b010;
		#2 b = 3'b111;
		$finish;
	end
/********************************************************************
 *                        MODULE IN TEST                            *
 *******************************************************************/
	top tops(a, b, c);
endmodule
